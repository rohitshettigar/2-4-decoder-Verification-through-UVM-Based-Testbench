interface deco_if ( input logic clk , reset ) ;
logic [1:0] in ;

logic [3:0] out ;

endinterface
