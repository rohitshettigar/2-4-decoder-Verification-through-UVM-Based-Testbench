class transaction ;
  bit [1:0] in ;
  bit [3:0] out ;
constraint in_c { in <4;}
endclass
